module weight_arrange(
  input i_clk,
  input i_rst_n,
  input [127:0] i_src_W_0,
  input [127:0] i_src_W_1,
  input [127:0] i_src_W_2,
  input [127:0] i_src_W_3,
  input [1:0] i_W_arrange,    
  input [1:0] i_W_arrange_index,
  output reg [31:0] o_W0,
  output reg [31:0] o_W1,
  output reg [31:0] o_W2,
  output reg [31:0] o_W3,
  output reg [31:0] o_W4,
  output reg [31:0] o_W5,
  output reg [31:0] o_W6,
  output reg [31:0] o_W7,
  output reg [31:0] o_W8,
  output reg [31:0] o_W9,
  output reg [31:0] o_W10,
  output reg [31:0] o_W11,
  output reg [31:0] o_W12,
  output reg [31:0] o_W13,
  output reg [31:0] o_W14,
  output reg [31:0] o_W15
);

  reg [1:0] W0_0, W0_1, W0_2, W0_3, W0_4, W0_5, W0_6, W0_7, W0_8, W0_9, W0_10, W0_11, W0_12, W0_13, W0_14, W0_15;
  reg [1:0] W1_0, W1_1, W1_2, W1_3, W1_4, W1_5, W1_6, W1_7, W1_8, W1_9, W1_10, W1_11, W1_12, W1_13, W1_14, W1_15;
  reg [1:0] W2_0, W2_1, W2_2, W2_3, W2_4, W2_5, W2_6, W2_7, W2_8, W2_9, W2_10, W2_11, W2_12, W2_13, W2_14, W2_15;
  reg [1:0] W3_0, W3_1, W3_2, W3_3, W3_4, W3_5, W3_6, W3_7, W3_8, W3_9, W3_10, W3_11, W3_12, W3_13, W3_14, W3_15;
  reg [1:0] W4_0, W4_1, W4_2, W4_3, W4_4, W4_5, W4_6, W4_7, W4_8, W4_9, W4_10, W4_11, W4_12, W4_13, W4_14, W4_15;
  reg [1:0] W5_0, W5_1, W5_2, W5_3, W5_4, W5_5, W5_6, W5_7, W5_8, W5_9, W5_10, W5_11, W5_12, W5_13, W5_14, W5_15;
  reg [1:0] W6_0, W6_1, W6_2, W6_3, W6_4, W6_5, W6_6, W6_7, W6_8, W6_9, W6_10, W6_11, W6_12, W6_13, W6_14, W6_15;
  reg [1:0] W7_0, W7_1, W7_2, W7_3, W7_4, W7_5, W7_6, W7_7, W7_8, W7_9, W7_10, W7_11, W7_12, W7_13, W7_14, W7_15;
  reg [1:0] W8_0, W8_1, W8_2, W8_3, W8_4, W8_5, W8_6, W8_7, W8_8, W8_9, W8_10, W8_11, W8_12, W8_13, W8_14, W8_15;
  reg [1:0] W9_0, W9_1, W9_2, W9_3, W9_4, W9_5, W9_6, W9_7, W9_8, W9_9, W9_10, W9_11, W9_12, W9_13, W9_14, W9_15;
  reg [1:0] W10_0, W10_1, W10_2, W10_3, W10_4, W10_5, W10_6, W10_7, W10_8, W10_9, W10_10, W10_11, W10_12, W10_13, W10_14, W10_15;
  reg [1:0] W11_0, W11_1, W11_2, W11_3, W11_4, W11_5, W11_6, W11_7, W11_8, W11_9, W11_10, W11_11, W11_12, W11_13, W11_14, W11_15;
  reg [1:0] W12_0, W12_1, W12_2, W12_3, W12_4, W12_5, W12_6, W12_7, W12_8, W12_9, W12_10, W12_11, W12_12, W12_13, W12_14, W12_15;
  reg [1:0] W13_0, W13_1, W13_2, W13_3, W13_4, W13_5, W13_6, W13_7, W13_8, W13_9, W13_10, W13_11, W13_12, W13_13, W13_14, W13_15;
  reg [1:0] W14_0, W14_1, W14_2, W14_3, W14_4, W14_5, W14_6, W14_7, W14_8, W14_9, W14_10, W14_11, W14_12, W14_13, W14_14, W14_15;
  reg [1:0] W15_0, W15_1, W15_2, W15_3, W15_4, W15_5, W15_6, W15_7, W15_8, W15_9, W15_10, W15_11, W15_12, W15_13, W15_14, W15_15;

  wire [31:0] W0_temp  = {W0_0, W1_0, W2_0, W3_0, W4_0, W5_0, W6_0, W7_0, W8_0, W9_0, W10_0, W11_0, W12_0, W13_0, W14_0, W15_0};
  wire [31:0] W1_temp  = {W0_1, W1_1, W2_1, W3_1, W4_1, W5_1, W6_1, W7_1, W8_1, W9_1, W10_1, W11_1, W12_1, W13_1, W14_1, W15_1};
  wire [31:0] W2_temp  = {W0_2, W1_2, W2_2, W3_2, W4_2, W5_2, W6_2, W7_2, W8_2, W9_2, W10_2, W11_2, W12_2, W13_2, W14_2, W15_2};
  wire [31:0] W3_temp  = {W0_3, W1_3, W2_3, W3_3, W4_3, W5_3, W6_3, W7_3, W8_3, W9_3, W10_3, W11_3, W12_3, W13_3, W14_3, W15_3};
  wire [31:0] W4_temp  = {W0_4, W1_4, W2_4, W3_4, W4_4, W5_4, W6_4, W7_4, W8_4, W9_4, W10_4, W11_4, W12_4, W13_4, W14_4, W15_4};
  wire [31:0] W5_temp  = {W0_5, W1_5, W2_5, W3_5, W4_5, W5_5, W6_5, W7_5, W8_5, W9_5, W10_5, W11_5, W12_5, W13_5, W14_5, W15_5};
  wire [31:0] W6_temp  = {W0_6, W1_6, W2_6, W3_6, W4_6, W5_6, W6_6, W7_6, W8_6, W9_6, W10_6, W11_6, W12_6, W13_6, W14_6, W15_6};
  wire [31:0] W7_temp  = {W0_7, W1_7, W2_7, W3_7, W4_7, W5_7, W6_7, W7_7, W8_7, W9_7, W10_7, W11_7, W12_7, W13_7, W14_7, W15_7};
  wire [31:0] W8_temp  = {W0_8, W1_8, W2_8, W3_8, W4_8, W5_8, W6_8, W7_8, W8_8, W9_8, W10_8, W11_8, W12_8, W13_8, W14_8, W15_8};
  wire [31:0] W9_temp  = {W0_9, W1_9, W2_9, W3_9, W4_9, W5_9, W6_9, W7_9, W8_9, W9_9, W10_9, W11_9, W12_9, W13_9, W14_9, W15_9};
  wire [31:0] W10_temp = {W0_10, W1_10, W2_10, W3_10, W4_10, W5_10, W6_10, W7_10, W8_10, W9_10, W10_10, W11_10, W12_10, W13_10, W14_10, W15_10};
  wire [31:0] W11_temp = {W0_11, W1_11, W2_11, W3_11, W4_11, W5_11, W6_11, W7_11, W8_11, W9_11, W10_11, W11_11, W12_11, W13_11, W14_11, W15_11};
  wire [31:0] W12_temp = {W0_12, W1_12, W2_12, W3_12, W4_12, W5_12, W6_12, W7_12, W8_12, W9_12, W10_12, W11_12, W12_12, W13_12, W14_12, W15_12};
  wire [31:0] W13_temp = {W0_13, W1_13, W2_13, W3_13, W4_13, W5_13, W6_13, W7_13, W8_13, W9_13, W10_13, W11_13, W12_13, W13_13, W14_13, W15_13};
  wire [31:0] W14_temp = {W0_14, W1_14, W2_14, W3_14, W4_14, W5_14, W6_14, W7_14, W8_14, W9_14, W10_14, W11_14, W12_14, W13_14, W14_14, W15_14};
  wire [31:0] W15_temp = {W0_15, W1_15, W2_15, W3_15, W4_15, W5_15, W6_15, W7_15, W8_15, W9_15, W10_15, W11_15, W12_15, W13_15, W14_15, W15_15};

  always@(posedge i_clk or negedge i_rst_n)begin
    if(!i_rst_n)begin
      o_W0  <= 32'd0;
      o_W1  <= 32'd0;
      o_W2  <= 32'd0;
      o_W3  <= 32'd0;
      o_W4  <= 32'd0;
      o_W5  <= 32'd0;
      o_W6  <= 32'd0;
      o_W7  <= 32'd0;
      o_W8  <= 32'd0;
      o_W9  <= 32'd0;
      o_W10 <= 32'd0;
      o_W11 <= 32'd0;
      o_W12 <= 32'd0;
      o_W13 <= 32'd0;
      o_W14 <= 32'd0;
      o_W15 <= 32'd0; 
    end else begin
      o_W0  <= W0_temp;
      o_W1  <= W1_temp;
      o_W2  <= W2_temp;
      o_W3  <= W3_temp;
      o_W4  <= W4_temp;
      o_W5  <= W5_temp;
      o_W6  <= W6_temp;
      o_W7  <= W7_temp;
      o_W8  <= W8_temp;
      o_W9  <= W9_temp;
      o_W10 <= W10_temp;
      o_W11 <= W11_temp;
      o_W12 <= W12_temp;
      o_W13 <= W13_temp;
      o_W14 <= W14_temp;
      o_W15 <= W15_temp;
    end
  end

  wire [127:0] W_for_now_8;
  assign W_for_now_8 = (i_W_arrange_index==2'd0) ? i_src_W_0 :
                       (i_W_arrange_index==2'd1) ? i_src_W_1 :
                       (i_W_arrange_index==2'd2) ? i_src_W_2 :
                       i_src_W_3;

  wire [127:0] W_for_now_4_0;
  assign W_for_now_4_0 = (i_W_arrange_index==2'd0) ? i_src_W_0 : i_src_W_2;
  wire [127:0] W_for_now_4_1;
  assign W_for_now_4_1 = (i_W_arrange_index==2'd0) ? i_src_W_1 : i_src_W_3;

  always@(*)begin
    case(i_W_arrange)
      2'b00:begin//22
        {W0_15, W0_14, W0_13, W0_12, W0_11, W0_10, W0_9, W0_8, W0_7, W0_6, W0_5, W0_4, W0_3, W0_2, W0_1, W0_0}                 = i_src_W_0[31:0];
        {W1_15, W1_14, W1_13, W1_12, W1_11, W1_10, W1_9, W1_8, W1_7, W1_6, W1_5, W1_4, W1_3, W1_2, W1_1, W1_0}                 = i_src_W_0[63:32];
        {W2_15, W2_14, W2_13, W2_12, W2_11, W2_10, W2_9, W2_8, W2_7, W2_6, W2_5, W2_4, W2_3, W2_2, W2_1, W2_0}                 = i_src_W_0[95:64];
        {W3_15, W3_14, W3_13, W3_12, W3_11, W3_10, W3_9, W3_8, W3_7, W3_6, W3_5, W3_4, W3_3, W3_2, W3_1, W3_0}                 = i_src_W_0[127:96];
        {W4_15, W4_14, W4_13, W4_12, W4_11, W4_10, W4_9, W4_8, W4_7, W4_6, W4_5, W4_4, W4_3, W4_2, W4_1, W4_0}                 = i_src_W_1[31:0];
        {W5_15, W5_14, W5_13, W5_12, W5_11, W5_10, W5_9, W5_8, W5_7, W5_6, W5_5, W5_4, W5_3, W5_2, W5_1, W5_0}                 = i_src_W_1[63:32];
        {W6_15, W6_14, W6_13, W6_12, W6_11, W6_10, W6_9, W6_8, W6_7, W6_6, W6_5, W6_4, W6_3, W6_2, W6_1, W6_0}                 = i_src_W_1[95:64];
        {W7_15, W7_14, W7_13, W7_12, W7_11, W7_10, W7_9, W7_8, W7_7, W7_6, W7_5, W7_4, W7_3, W7_2, W7_1, W7_0}                 = i_src_W_1[127:96];
        {W8_15, W8_14, W8_13, W8_12, W8_11, W8_10, W8_9, W8_8, W8_7, W8_6, W8_5, W8_4, W8_3, W8_2, W8_1, W8_0}                 = i_src_W_2[31:0];
        {W9_15, W9_14, W9_13, W9_12, W9_11, W9_10, W9_9, W9_8, W9_7, W9_6, W9_5, W9_4, W9_3, W9_2, W9_1, W9_0}                 = i_src_W_2[63:32];
        {W10_15, W10_14, W10_13, W10_12, W10_11, W10_10, W10_9, W10_8, W10_7, W10_6, W10_5, W10_4, W10_3, W10_2, W10_1, W10_0} = i_src_W_2[95:64];
        {W11_15, W11_14, W11_13, W11_12, W11_11, W11_10, W11_9, W11_8, W11_7, W11_6, W11_5, W11_4, W11_3, W11_2, W11_1, W11_0} = i_src_W_2[127:96];
        {W12_15, W12_14, W12_13, W12_12, W12_11, W12_10, W12_9, W12_8, W12_7, W12_6, W12_5, W12_4, W12_3, W12_2, W12_1, W12_0} = i_src_W_3[31:0];
        {W13_15, W13_14, W13_13, W13_12, W13_11, W13_10, W13_9, W13_8, W13_7, W13_6, W13_5, W13_4, W13_3, W13_2, W13_1, W13_0} = i_src_W_3[63:32];
        {W14_15, W14_14, W14_13, W14_12, W14_11, W14_10, W14_9, W14_8, W14_7, W14_6, W14_5, W14_4, W14_3, W14_2, W14_1, W14_0} = i_src_W_3[95:64];
        {W15_15, W15_14, W15_13, W15_12, W15_11, W15_10, W15_9, W15_8, W15_7, W15_6, W15_5, W15_4, W15_3, W15_2, W15_1, W15_0} = i_src_W_3[127:96];
      end
      2'b01:begin//42
        {W0_14, W0_12, W0_10, W0_8, W0_15, W0_13, W0_11, W0_9, W0_6, W0_4, W0_2, W0_0, W0_7, W0_5, W0_3, W0_1}                 = {W_for_now_4_0[15:8], W_for_now_4_0[15:8], W_for_now_4_0[7:0], W_for_now_4_0[7:0]};
        {W1_14, W1_12, W1_10, W1_8, W1_15, W1_13, W1_11, W1_9, W1_6, W1_4, W1_2, W1_0, W1_7, W1_5, W1_3, W1_1}                 = {W_for_now_4_0[31:24], W_for_now_4_0[31:24], W_for_now_4_0[23:16], W_for_now_4_0[23:16]};
        {W2_14, W2_12, W2_10, W2_8, W2_15, W2_13, W2_11, W2_9, W2_6, W2_4, W2_2, W2_0, W2_7, W2_5, W2_3, W2_1}                 = {W_for_now_4_0[47:40], W_for_now_4_0[47:40], W_for_now_4_0[39:32], W_for_now_4_0[39:32]};
        {W3_14, W3_12, W3_10, W3_8, W3_15, W3_13, W3_11, W3_9, W3_6, W3_4, W3_2, W3_0, W3_7, W3_5, W3_3, W3_1}                 = {W_for_now_4_0[63:56], W_for_now_4_0[63:56], W_for_now_4_0[55:48], W_for_now_4_0[55:48]};
        {W4_14, W4_12, W4_10, W4_8, W4_15, W4_13, W4_11, W4_9, W4_6, W4_4, W4_2, W4_0, W4_7, W4_5, W4_3, W4_1}                 = {W_for_now_4_0[79:72], W_for_now_4_0[79:72], W_for_now_4_0[71:64], W_for_now_4_0[71:64]};
        {W5_14, W5_12, W5_10, W5_8, W5_15, W5_13, W5_11, W5_9, W5_6, W5_4, W5_2, W5_0, W5_7, W5_5, W5_3, W5_1}                 = {W_for_now_4_0[95:88], W_for_now_4_0[95:88], W_for_now_4_0[87:80], W_for_now_4_0[87:80]};
        {W6_14, W6_12, W6_10, W6_8, W6_15, W6_13, W6_11, W6_9, W6_6, W6_4, W6_2, W6_0, W6_7, W6_5, W6_3, W6_1}                 = {W_for_now_4_0[111:104], W_for_now_4_0[111:104], W_for_now_4_0[103:96], W_for_now_4_0[103:96]};
        {W7_14, W7_12, W7_10, W7_8, W7_15, W7_13, W7_11, W7_9, W7_6, W7_4, W7_2, W7_0, W7_7, W7_5, W7_3, W7_1}                 = {W_for_now_4_0[127:120], W_for_now_4_0[127:120], W_for_now_4_0[119:112], W_for_now_4_0[119:112]};
        {W8_14, W8_12, W8_10, W8_8, W8_15, W8_13, W8_11, W8_9, W8_6, W8_4, W8_2, W8_0, W8_7, W8_5, W8_3, W8_1}                 = {W_for_now_4_1[15:8], W_for_now_4_1[15:8], W_for_now_4_1[7:0], W_for_now_4_1[7:0]};
        {W9_14, W9_12, W9_10, W9_8, W9_15, W9_13, W9_11, W9_9, W9_6, W9_4, W9_2, W9_0, W9_7, W9_5, W9_3, W9_1}                 = {W_for_now_4_1[31:24], W_for_now_4_1[31:24], W_for_now_4_1[23:16], W_for_now_4_1[23:16]};
        {W10_14, W10_12, W10_10, W10_8, W10_15, W10_13, W10_11, W10_9, W10_6, W10_4, W10_2, W10_0, W10_7, W10_5, W10_3, W10_1} = {W_for_now_4_1[47:40], W_for_now_4_1[47:40], W_for_now_4_1[39:32], W_for_now_4_1[39:32]};
        {W11_14, W11_12, W11_10, W11_8, W11_15, W11_13, W11_11, W11_9, W11_6, W11_4, W11_2, W11_0, W11_7, W11_5, W11_3, W11_1} = {W_for_now_4_1[63:56], W_for_now_4_1[63:56], W_for_now_4_1[55:48], W_for_now_4_1[55:48]};
        {W12_14, W12_12, W12_10, W12_8, W12_15, W12_13, W12_11, W12_9, W12_6, W12_4, W12_2, W12_0, W12_7, W12_5, W12_3, W12_1} = {W_for_now_4_1[79:72], W_for_now_4_1[79:72], W_for_now_4_1[71:64], W_for_now_4_1[71:64]};
        {W13_14, W13_12, W13_10, W13_8, W13_15, W13_13, W13_11, W13_9, W13_6, W13_4, W13_2, W13_0, W13_7, W13_5, W13_3, W13_1} = {W_for_now_4_1[95:88], W_for_now_4_1[95:88], W_for_now_4_1[87:80], W_for_now_4_1[87:80]};
        {W14_14, W14_12, W14_10, W14_8, W14_15, W14_13, W14_11, W14_9, W14_6, W14_4, W14_2, W14_0, W14_7, W14_5, W14_3, W14_1} = {W_for_now_4_1[111:104], W_for_now_4_1[111:104], W_for_now_4_1[103:96], W_for_now_4_1[103:96]};
        {W15_14, W15_12, W15_10, W15_8, W15_15, W15_13, W15_11, W15_9, W15_6, W15_4, W15_2, W15_0, W15_7, W15_5, W15_3, W15_1} = {W_for_now_4_1[127:120], W_for_now_4_1[127:120], W_for_now_4_1[119:112], W_for_now_4_1[119:112]};
      end
      2'b10:begin//44
        {W0_14, W0_10, W0_12, W0_8, W0_15, W0_11, W0_13, W0_9, W0_6, W0_2, W0_4, W0_0, W0_7, W0_3, W0_5, W0_1}                 = {W_for_now_4_0[15:8], W_for_now_4_0[15:8], W_for_now_4_0[7:0], W_for_now_4_0[7:0]};
        {W1_14, W1_10, W1_12, W1_8, W1_15, W1_11, W1_13, W1_9, W1_6, W1_2, W1_4, W1_0, W1_7, W1_3, W1_5, W1_1}                 = {W_for_now_4_0[31:24], W_for_now_4_0[31:24], W_for_now_4_0[23:16], W_for_now_4_0[23:16]};
        {W2_14, W2_10, W2_12, W2_8, W2_15, W2_11, W2_13, W2_9, W2_6, W2_2, W2_4, W2_0, W2_7, W2_3, W2_5, W2_1}                 = {W_for_now_4_0[47:40], W_for_now_4_0[47:40], W_for_now_4_0[39:32], W_for_now_4_0[39:32]};
        {W3_14, W3_10, W3_12, W3_8, W3_15, W3_11, W3_13, W3_9, W3_6, W3_2, W3_4, W3_0, W3_7, W3_3, W3_5, W3_1}                 = {W_for_now_4_0[63:56], W_for_now_4_0[63:56], W_for_now_4_0[55:48], W_for_now_4_0[55:48]};
        {W4_14, W4_10, W4_12, W4_8, W4_15, W4_11, W4_13, W4_9, W4_6, W4_2, W4_4, W4_0, W4_7, W4_3, W4_5, W4_1}                 = {W_for_now_4_0[79:72], W_for_now_4_0[79:72], W_for_now_4_0[71:64], W_for_now_4_0[71:64]};
        {W5_14, W5_10, W5_12, W5_8, W5_15, W5_11, W5_13, W5_9, W5_6, W5_2, W5_4, W5_0, W5_7, W5_3, W5_5, W5_1}                 = {W_for_now_4_0[95:88], W_for_now_4_0[95:88], W_for_now_4_0[87:80], W_for_now_4_0[87:80]};
        {W6_14, W6_10, W6_12, W6_8, W6_15, W6_11, W6_13, W6_9, W6_6, W6_2, W6_4, W6_0, W6_7, W6_3, W6_5, W6_1}                 = {W_for_now_4_0[111:104], W_for_now_4_0[111:104], W_for_now_4_0[103:96], W_for_now_4_0[103:96]};
        {W7_14, W7_10, W7_12, W7_8, W7_15, W7_11, W7_13, W7_9, W7_6, W7_2, W7_4, W7_0, W7_7, W7_3, W7_5, W7_1}                 = {W_for_now_4_0[127:120], W_for_now_4_0[127:120], W_for_now_4_0[119:112], W_for_now_4_0[119:112]};
        {W8_14, W8_10, W8_12, W8_8, W8_15, W8_11, W8_13, W8_9, W8_6, W8_2, W8_4, W8_0, W8_7, W8_3, W8_5, W8_1}                 = {W_for_now_4_1[15:8], W_for_now_4_1[15:8], W_for_now_4_1[7:0], W_for_now_4_1[7:0]};
        {W9_14, W9_10, W9_12, W9_8, W9_15, W9_11, W9_13, W9_9, W9_6, W9_2, W9_4, W9_0, W9_7, W9_3, W9_5, W9_1}                 = {W_for_now_4_1[31:24], W_for_now_4_1[31:24], W_for_now_4_1[23:16], W_for_now_4_1[23:16]};
        {W10_14, W10_10, W10_12, W10_8, W10_15, W10_11, W10_13, W10_9, W10_6, W10_2, W10_4, W10_0, W10_7, W10_3, W10_5, W10_1} = {W_for_now_4_1[47:40], W_for_now_4_1[47:40], W_for_now_4_1[39:32], W_for_now_4_1[39:32]};
        {W11_14, W11_10, W11_12, W11_8, W11_15, W11_11, W11_13, W11_9, W11_6, W11_2, W11_4, W11_0, W11_7, W11_3, W11_5, W11_1} = {W_for_now_4_1[63:56], W_for_now_4_1[63:56], W_for_now_4_1[55:48], W_for_now_4_1[55:48]};
        {W12_14, W12_10, W12_12, W12_8, W12_15, W12_11, W12_13, W12_9, W12_6, W12_2, W12_4, W12_0, W12_7, W12_3, W12_5, W12_1} = {W_for_now_4_1[79:72], W_for_now_4_1[79:72], W_for_now_4_1[71:64], W_for_now_4_1[71:64]};
        {W13_14, W13_10, W13_12, W13_8, W13_15, W13_11, W13_13, W13_9, W13_6, W13_2, W13_4, W13_0, W13_7, W13_3, W13_5, W13_1} = {W_for_now_4_1[95:88], W_for_now_4_1[95:88], W_for_now_4_1[87:80], W_for_now_4_1[87:80]};
        {W14_14, W14_10, W14_12, W14_8, W14_15, W14_11, W14_13, W14_9, W14_6, W14_2, W14_4, W14_0, W14_7, W14_3, W14_5, W14_1} = {W_for_now_4_1[111:104], W_for_now_4_1[111:104], W_for_now_4_1[103:96], W_for_now_4_1[103:96]};
        {W15_14, W15_10, W15_12, W15_8, W15_15, W15_11, W15_13, W15_9, W15_6, W15_2, W15_4, W15_0, W15_7, W15_3, W15_5, W15_1} = {W_for_now_4_1[127:120], W_for_now_4_1[127:120], W_for_now_4_1[119:112], W_for_now_4_1[119:112]};
      end
      default:begin//88 84 82
        {W0_12, W0_8, W0_4, W0_0, W0_13, W0_9, W0_5, W0_1, W0_14, W0_10, W0_6, W0_2, W0_15, W0_11, W0_7, W0_3}                 = {W_for_now_8[7:0], W_for_now_8[7:0], W_for_now_8[7:0], W_for_now_8[7:0]};      
        {W1_12, W1_8, W1_4, W1_0, W1_13, W1_9, W1_5, W1_1, W1_14, W1_10, W1_6, W1_2, W1_15, W1_11, W1_7, W1_3}                 = {W_for_now_8[15:8], W_for_now_8[15:8], W_for_now_8[15:8], W_for_now_8[15:8]};
        {W2_12, W2_8, W2_4, W2_0, W2_13, W2_9, W2_5, W2_1, W2_14, W2_10, W2_6, W2_2, W2_15, W2_11, W2_7, W2_3}                 = {W_for_now_8[23:16], W_for_now_8[23:16], W_for_now_8[23:16], W_for_now_8[23:16]};
        {W3_12, W3_8, W3_4, W3_0, W3_13, W3_9, W3_5, W3_1, W3_14, W3_10, W3_6, W3_2, W3_15, W3_11, W3_7, W3_3}                 = {W_for_now_8[31:24], W_for_now_8[31:24], W_for_now_8[31:24], W_for_now_8[31:24]};
        {W4_12, W4_8, W4_4, W4_0, W4_13, W4_9, W4_5, W4_1, W4_14, W4_10, W4_6, W4_2, W4_15, W4_11, W4_7, W4_3}                 = {W_for_now_8[39:32], W_for_now_8[39:32], W_for_now_8[39:32], W_for_now_8[39:32]};
        {W5_12, W5_8, W5_4, W5_0, W5_13, W5_9, W5_5, W5_1, W5_14, W5_10, W5_6, W5_2, W5_15, W5_11, W5_7, W5_3}                 = {W_for_now_8[47:40], W_for_now_8[47:40], W_for_now_8[47:40], W_for_now_8[47:40]};
        {W6_12, W6_8, W6_4, W6_0, W6_13, W6_9, W6_5, W6_1, W6_14, W6_10, W6_6, W6_2, W6_15, W6_11, W6_7, W6_3}                 = {W_for_now_8[55:48], W_for_now_8[55:48], W_for_now_8[55:48], W_for_now_8[55:48]};
        {W7_12, W7_8, W7_4, W7_0, W7_13, W7_9, W7_5, W7_1, W7_14, W7_10, W7_6, W7_2, W7_15, W7_11, W7_7, W7_3}                 = {W_for_now_8[63:56], W_for_now_8[63:56], W_for_now_8[63:56], W_for_now_8[63:56]};
        {W8_12, W8_8, W8_4, W8_0, W8_13, W8_9, W8_5, W8_1, W8_14, W8_10, W8_6, W8_2, W8_15, W8_11, W8_7, W8_3}                 = {W_for_now_8[71:64], W_for_now_8[71:64], W_for_now_8[71:64], W_for_now_8[71:64]};
        {W9_12, W9_8, W9_4, W9_0, W9_13, W9_9, W9_5, W9_1, W9_14, W9_10, W9_6, W9_2, W9_15, W9_11, W9_7, W9_3}                 = {W_for_now_8[79:72], W_for_now_8[79:72], W_for_now_8[79:72], W_for_now_8[79:72]};
        {W10_12, W10_8, W10_4, W10_0, W10_13, W10_9, W10_5, W10_1, W10_14, W10_10, W10_6, W10_2, W10_15, W10_11, W10_7, W10_3} = {W_for_now_8[87:80], W_for_now_8[87:80], W_for_now_8[87:80], W_for_now_8[87:80]};
        {W11_12, W11_8, W11_4, W11_0, W11_13, W11_9, W11_5, W11_1, W11_14, W11_10, W11_6, W11_2, W11_15, W11_11, W11_7, W11_3} = {W_for_now_8[95:88], W_for_now_8[95:88], W_for_now_8[95:88], W_for_now_8[95:88]};
        {W12_12, W12_8, W12_4, W12_0, W12_13, W12_9, W12_5, W12_1, W12_14, W12_10, W12_6, W12_2, W12_15, W12_11, W12_7, W12_3} = {W_for_now_8[103:96], W_for_now_8[103:96], W_for_now_8[103:96], W_for_now_8[103:96]};
        {W13_12, W13_8, W13_4, W13_0, W13_13, W13_9, W13_5, W13_1, W13_14, W13_10, W13_6, W13_2, W13_15, W13_11, W13_7, W13_3} = {W_for_now_8[111:104], W_for_now_8[111:104], W_for_now_8[111:104], W_for_now_8[111:104]};
        {W14_12, W14_8, W14_4, W14_0, W14_13, W14_9, W14_5, W14_1, W14_14, W14_10, W14_6, W14_2, W14_15, W14_11, W14_7, W14_3} = {W_for_now_8[119:112], W_for_now_8[119:112], W_for_now_8[119:112], W_for_now_8[119:112]};
        {W15_12, W15_8, W15_4, W15_0, W15_13, W15_9, W15_5, W15_1, W15_14, W15_10, W15_6, W15_2, W15_15, W15_11, W15_7, W15_3} = {W_for_now_8[127:120], W_for_now_8[127:120], W_for_now_8[127:120], W_for_now_8[127:120]};
      end
    endcase
  end

endmodule